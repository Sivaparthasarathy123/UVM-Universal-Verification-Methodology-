// ASYNCHRONOUS FIFO - UVM PARAMETER PACKAGE

`ifndef ASYNC_FIFO_PKG_SV
`define ASYNC_FIFO_PKG_SV

package async_fifo_pkg;
  parameter DEPTH = 8;
  parameter WIDTH = 8;
endpackage

`endif
