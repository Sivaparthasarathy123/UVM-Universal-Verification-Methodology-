// SYNCHRONOUS FIFO - UVM PARAMETER PACKAGE
`ifndef SYNC_FIFO_PKG_SV
`define SYNC_FIFO_PKG_SV

package sync_fifo_pkg;
  parameter DEPTH = 16;
  parameter WIDTH = 16;
endpackage

`endif
